`ifndef DEFINES_VH
`define DEFINES_VH

`timescale 1ns/1ps

`endif