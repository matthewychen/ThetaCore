module CU_SV();

endmodule