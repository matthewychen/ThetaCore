module CU_decrypt(
    input [31:0] CU_in,
    output [4:0] module_sel,
    output [31:0] CU_to_ALU,

);//deprecate. ALU should be instantiated in CU

endmodule