module SRAM(
    input [7:0] addr,
    input [31:0] datain,
    output [31:0] dataout,
    output f_ready
);



endmodule