module memfetch(
    //templated
    input soc_clk,
    input reset,
    input CU_ready
    //need to retrieve from and write data to SRAM.
);

endmodule