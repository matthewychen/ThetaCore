module ALU_top(
    input sysclk,
    input [31:0] ALU_dat1,
    input [31:0] ALU_dat2,
    input [7:0] ALU_op,

    //flags
    output ALU_underflow,
    output ALU_overflow,
    output ALU_out
    );

    

endmodule