module CU_MEM(
    
);

// need to edit and pass signals back upwards to interface with MMU

endmodule