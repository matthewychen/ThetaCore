module CU_MEM(
    
);

endmodule