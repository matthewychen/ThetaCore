module ControlUnit(

);

CU_decrpyt CU_decrypt_inst(
    .CU_out(CU_out)
);

endmodule